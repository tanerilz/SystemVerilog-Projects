package env_package;
   import agent_package::*;
   import uvm_pkg::*;
`include "uvm_macros.svh"
`include "scoreboard.svh"
`include "env_cfg.svh"
`include "env.svh"
endpackage // Environment_package
   