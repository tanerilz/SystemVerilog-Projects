package Environment_package;
   import agent_package::*;
   
`include "scoreboard.svh"
`include "environment.svh"
endpackage // Environment_package
   