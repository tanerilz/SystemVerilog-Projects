interface iface(input logic clock, reset);
   bit s1,s2;
   bit light;
   bit full,empty;
endinterface
 	