package test_package;
   import environment_package::*;
   import uvm_pkg::*;
   import agent_package::*;
`include "test.svh"

endpackage // test_package
   