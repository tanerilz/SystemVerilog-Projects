package environment_package;
   import agent_package::*;
   import uvm_pkg::*;
`include "uvm_macros.svh"
`include "scoreboard.svh"
`include "environment_cfg.svh"
`include "environment.svh"
endpackage // Environment_package
   