class Transaction;
   rand logic  write_req,read_req;
   rand logic [7:0] write_data;
   logic [7:0] read_data;
   logic       FULL,EMP;
endclass:Transaction
