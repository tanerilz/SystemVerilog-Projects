package agent_package;
`include "transaction.svh"
`include "generator.svh"
`include "driver.svh"
`include "monitor.svh"
`include "agent.svh"
endpackage // agent_package
   