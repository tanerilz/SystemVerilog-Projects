package agent_package;
 import uvm_pkg::*;
`include "uvm_macros.svh"
`include "transaction.svh"
`include "agent_cfg.svh"
`include "sequence.svh"
`include "sequencer.svh"
`include "driver.svh"
`include "monitor.svh"
`include "agent.svh"
endpackage // agent_package
   